import uvm_pkg::*;

`include "ialu_base_seq_item_pkg.svh"
`include "ialu_sum1_seq_item_pkg.svh"

`include "ialu_base_sequencer_config_pkg.svh"
`include "ialu_base_sequencer_pkg.svh"
`include "ialu_sum1_sequencer_config_pkg.svh"
`include "ialu_sum1_sequencer_pkg.svh"

`include "ialu_base_sequence_pkg.svh"
`include "ialu_sum1_sequence_pkg.svh"

`include "ialu_base_driver_pkg.svh"
`include "ialu_sum1_driver_pkg.svh"

`include "ialu_base_monitor_pkg.svh"
`include "ialu_sum1_monitor_pkg.svh"

`include "ialu_scoreboard_config_pkg.svh"
`include "ialu_scoreboard_pkg.svh"

`include "ialu_base_agent_config_pkg.svh"
`include "ialu_base_agent_pkg.svh"
`include "ialu_sum1_agent_config_pkg.svh"
`include "ialu_sum1_agent_pkg.svh"

`include "ialu_env_config_pkg.svh"
`include "ialu_env_pkg.svh"

`include "ialu_base_test_pkg.svh"
`include "ialu_full_test_pkg.svh"
