`ifndef IALU_BASE_SEQUENCER_CONFIG
`define IALU_BASE_SEQUENCER_CONFIG

virtual class ialu_base_sequencer_config extends uvm_object;
  // ---------------------------------------------------------------------------
  // Members
  // ---------------------------------------------------------------------------
  //
  // ---------------------------------------------------------------------------
  // Class Methods
  // ---------------------------------------------------------------------------
  //
  // ---------------------------------------------------------------------------
  //                                                                 UVM Methods
  // ---------------------------------------------------------------------------
  //
  extern function new (string name = "ialu_base_sequencer_config");


endclass : ialu_base_sequencer_config