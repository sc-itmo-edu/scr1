
class ialu_sum1_sequencer_config extends ialu_base_sequencer_config;
  `uvm_object_utils(ialu_sum1_sequencer_config)
  // ---------------------------------------------------------------------------
  // Members
  // ---------------------------------------------------------------------------
  //
  // ---------------------------------------------------------------------------
  // Class Methods
  // ---------------------------------------------------------------------------
  //
  // ---------------------------------------------------------------------------
  //                                                                 UVM Methods
  // ---------------------------------------------------------------------------
  //
  extern function new (string name = "ialu_sum1_sequencer_config");


endclass : ialu_sum1_sequencer_config