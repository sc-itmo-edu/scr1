`include "ialu_tb_pkg.svh"

`include "scr1_pipe_ialu.sv"

`include "ialu_sum1_if.sv"
`include "ialu_tb_lib.sv"
`include "ialu_wrapper.sv"
`include "ialu_tb_top.sv"